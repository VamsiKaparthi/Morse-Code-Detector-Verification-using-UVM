package pkg;
	`include "uvm_macros.svh"
	import uvm_pkg::*;
	`include "mor_seq_item.sv";
endpackage
