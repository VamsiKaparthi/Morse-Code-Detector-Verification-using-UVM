parameter N = 1;
