package pkg;
	`include "uvm_macros.svh"
	import uvm_pkg::*;
	`include "define.svh";
	`include "mor_seq_item.sv";
	`include "mor_sequence.sv";
	`include "mor_sequencer.sv";
	`include "mor_driver.sv";
	`include "mor_monitor.sv";
	`include "mor_agent.sv";
endpackage
